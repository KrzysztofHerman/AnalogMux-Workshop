** sch_path: /home/herman/tmp/ts_pr_May2024/design_data/xschem/transmission_gate_tb_On-Off-time.sch
**.subckt transmission_gate_tb_On-Off-time
Vpow Vdd GND 1.2
Vp Vdd net1 0
.save i(vp)
Vin V_in GND dc=0 ac=1 pulse(0 1.2 25n 1p 1p 105n 110n)
Ven en_p GND pulse(0 1.2 50n 1p 1p 50n 100n)
C1 V_out GND 1p m=1
Ven1 en_n GND pulse(0 1.2 0 1p 1p 50n 100n)
x1 net1 en_n V_in V_out en_p GND transmission_gate
R1 V_out GND 10k m=1
**** begin user architecture code

.lib cornerMOSlv.lib mos_tt
.lib cornerRES.lib res_typ



.param temp=27
.control
save all
tran 10p 150n
meas tran turn-On TRIG v(en_p) VAL=0.6 RISE=1 TARG v(v_out) VAL=1.1 RISE=1
meas tran turn-OFF TRIG v(en_p) VAL=0.6 FALL=1 TARG v(v_out) VAL=0.1 FALL=1
write tran_ton-off.raw
set hcopydevtype=svg
set color0=white
set color1=black
set color2=red
set color3=blue
set color4=green
hardcopy turn-on-off1.svg en_p v_out title 'Turn On/Off time' xlabel 'time' ylabel 'voltage'
hardcopy turn-on-off2.svg v_in v_out title 'Turn On/Off time' xlabel 'time' ylabel 'voltage'

.endc


**** end user architecture code
**.ends

* expanding   symbol:  transmission_gate.sym # of pins=6
** sym_path: /home/herman/tmp/ts_pr_May2024/design_data/xschem/transmission_gate.sym
** sch_path: /home/herman/tmp/ts_pr_May2024/design_data/xschem/transmission_gate.sch
.subckt transmission_gate vdd en_n inout_1 inout_2 en_p vss
*.iopin inout_1
*.iopin inout_2
*.ipin en_p
*.iopin vdd
*.iopin vss
*.ipin en_n
XM1 inout_2 en_p inout_1 net1 sg13_lv_nmos w=200.0u l=0.130u ng=20 m=1
XM2 inout_1 en_n inout_2 net2 sg13_lv_pmos w=200.0u l=0.130u ng=20 m=1
XR1 net2 vdd ntap1
XR2 net1 vss ptap1
.ends

.GLOBAL GND
.end
