** sch_path: /home/herman/tmp/ts_pr_May2024/design_data/xschem/transmission_gate_tb_noise.sch
**.subckt transmission_gate_tb_noise
Vpow Vdd GND 1.2
Vp Vdd net1 0
.save i(vp)
Vin V_in GND dc 0 ac 1
Ven en_p GND 1.2
Ven1 en_n GND 0
x1 net1 en_n V_in V_out en_p GND transmission_gate
R1 V_out GND 50 m=1
**** begin user architecture code

.lib cornerMOSlv.lib mos_tt
.lib cornerRES.lib res_typ



.param temp=27
.control
save all
noise V(V_out) Vin dec 1001 10 10G
setplot noise1
set hcopydevtype=svg
set color0=white
set color1=black
set color2=red
set color3=blue
set color4=green
hardcopy noise1.svg onoise_spectrum  title 'Output noise spectrum' xlabel 'frequency' ylabel 'Vout' xlog
setplot noise2
print onoise_total
.endc


**** end user architecture code
**.ends

* expanding   symbol:  transmission_gate.sym # of pins=6
** sym_path: /home/herman/tmp/ts_pr_May2024/design_data/xschem/transmission_gate.sym
** sch_path: /home/herman/tmp/ts_pr_May2024/design_data/xschem/transmission_gate.sch
.subckt transmission_gate vdd en_n inout_1 inout_2 en_p vss
*.iopin inout_1
*.iopin inout_2
*.ipin en_p
*.iopin vdd
*.iopin vss
*.ipin en_n
XM1 inout_2 en_p inout_1 net1 sg13_lv_nmos w=200.0u l=0.130u ng=20 m=1
XM2 inout_1 en_n inout_2 net2 sg13_lv_pmos w=200.0u l=0.130u ng=20 m=1
XR1 net2 vdd ntap1
XR2 net1 vss ptap1
.ends

.GLOBAL GND
.end
