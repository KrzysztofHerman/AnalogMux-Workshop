module multiplexer(
  
  input [7:0] analog_i,
  output analog_o,
  input [15:0] ctrl
);

endmodule
