** sch_path: /home/herman/tmp/ts_pr_May2024/design_data/xschem/transmission_gate_tb_Ileak.sch
**.subckt transmission_gate_tb_Ileak
Vpow Vdd GND 1.2
Vp Vdd net3 0
.save i(vp)
Vin V_in GND 0
Ven en_p GND 0
Ven1 en_n GND 1.2
x1 net3 en_n net2 net1 en_p GND transmission_gate
Vout V_out1 GND 1.2
Vp1 V_out1 net1 0
.save i(vp1)
Vp2 net2 V_in 0
.save i(vp2)
Vp3 Vdd net5 0
.save i(vp3)
x2 net5 en_p net4 V_out1 en_n GND transmission_gate
Vp5 net6 net4 0
.save i(vp5)
Vin1 net6 GND 1.2
**** begin user architecture code

.lib cornerMOSlv.lib mos_tt
.lib cornerRES.lib res_typ



.param temp=27
.control
save all
op
echo Off state leakage currents
echo output current
print I(Vp1)
echo input current
print I(Vp2)
echo on state leakage current
print I(Vp5)
write op_Ileak.raw
.endc


**** end user architecture code
**.ends

* expanding   symbol:  transmission_gate.sym # of pins=6
** sym_path: /home/herman/tmp/ts_pr_May2024/design_data/xschem/transmission_gate.sym
** sch_path: /home/herman/tmp/ts_pr_May2024/design_data/xschem/transmission_gate.sch
.subckt transmission_gate vdd en_n inout_1 inout_2 en_p vss
*.iopin inout_1
*.iopin inout_2
*.ipin en_p
*.iopin vdd
*.iopin vss
*.ipin en_n
XM1 inout_2 en_p inout_1 net1 sg13_lv_nmos w=200.0u l=0.130u ng=20 m=1
XM2 inout_1 en_n inout_2 net2 sg13_lv_pmos w=200.0u l=0.130u ng=20 m=1
XR1 net2 vdd ntap1
XR2 net1 vss ptap1
.ends

.GLOBAL GND
.end
