module bondpad_70x70 ();
endmodule
