** sch_path: /home/herman/tmp/ts_pr_May2024/design_data/xschem/transmission_gate_tb_Cinject.sch
**.subckt transmission_gate_tb_Cinject
Vpow Vdd GND 1.2
Vp Vdd net1 0
.save i(vp)
Vin V_in GND 1
Ven en_p GND pulse(0 1.2 50n 1p 1p 50n 100n)
C1 V_out GND 1p m=1
Ven1 en_n GND pulse(0 1.2 0 1p 1p 50n 100n)
x1 net1 en_n GND V_out en_p GND transmission_gate
**** begin user architecture code

.lib cornerMOSlv.lib mos_tt
.lib cornerRES.lib res_typ



.param temp=27
.control
save all
tran 10p 150n
write tran_cinject.raw
set hcopydevtype=svg
set color0=white
set color1=black
set color2=red
set color3=blue
set color4=green
hardcopy cinject1.svg v_out  title 'Output voltage' xlabel 'time' ylabel 'voltage'
hardcopy cinject2.svg en_p   title 'Control signal' xlabel 'time' ylabel 'voltage'

.endc


**** end user architecture code
**.ends

* expanding   symbol:  transmission_gate.sym # of pins=6
** sym_path: /home/herman/tmp/ts_pr_May2024/design_data/xschem/transmission_gate.sym
** sch_path: /home/herman/tmp/ts_pr_May2024/design_data/xschem/transmission_gate.sch
.subckt transmission_gate vdd en_n inout_1 inout_2 en_p vss
*.iopin inout_1
*.iopin inout_2
*.ipin en_p
*.iopin vdd
*.iopin vss
*.ipin en_n
XM1 inout_2 en_p inout_1 net1 sg13_lv_nmos w=200.0u l=0.130u ng=20 m=1
XM2 inout_1 en_n inout_2 net2 sg13_lv_pmos w=200.0u l=0.130u ng=20 m=1
XR1 net2 vdd ntap1
XR2 net1 vss ptap1
.ends

.GLOBAL GND
.end
